module test (a, ctrl, o);
  input a, ctrl;
  output o;
  pmos (o, a, ctrl);
endmodule
