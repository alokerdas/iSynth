module test (a, ctrl, o);
  input a, ctrl;
  output o;
  rpmos (o, a, ctrl);
endmodule
