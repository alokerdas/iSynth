module test (a, ctrl, o);
  input a, ctrl;
  output o;
  notif1 (o, a, ctrl);
endmodule
