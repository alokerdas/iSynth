module test (a, b, o);
  input [1:0] a, b;
  output [3:0]o;
  assign o = a * b;
endmodule
