module test (a, ctrl, o);
  input a, ctrl;
  output o;
  nmos (o, a, ctrl);
endmodule
