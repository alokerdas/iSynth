module test (a, ctrl, o);
  input a, ctrl;
  output o;
  tranif1 (a, o, ctrl);
endmodule
