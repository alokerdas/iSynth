module test (a, ctrl, o);
  input a, ctrl;
  output o;
  tranif0 (a, o, ctrl);
endmodule
