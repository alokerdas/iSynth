module test (a, o);
  input a;
  output o;
  tran (a, o);
endmodule
