module test (o);
  integer a;
  output o;
  assign o = abs(a);
endmodule
