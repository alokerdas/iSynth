module test (a, ctrl, o);
  input a, ctrl;
  output o;
  rtranif1 (a, o, ctrl);
endmodule
