module test (a, o);
  input a;
  output o;
  rtran (a, o);
endmodule
