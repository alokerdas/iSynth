module test (a, ctrl, o);
  input a, ctrl;
  output o;
  rnmos (o, a, ctrl);
endmodule
