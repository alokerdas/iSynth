module test (o, a, b);
  input a, b;
  output o;
  assign o = a >= b;
endmodule
