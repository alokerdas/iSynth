module test (a, ctrl, o);
  input a, ctrl;
  output o;
  notif0 (o, a, ctrl);
endmodule
