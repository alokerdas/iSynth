module test (a, b, o);
  input [1:0] a;
  input b;
  output [2:0] o;
  assign o = a * b;
endmodule
