module test (a, ctrl, o);
  input a, ctrl;
  output o;
  rtranif0 (a, o, ctrl);
endmodule
